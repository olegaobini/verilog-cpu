
module DmemReg();
    input logic [7:0] D_addr
endmodule